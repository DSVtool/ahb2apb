// File name: 			bridge_macros.sv
// Creator name: 		Dimitrije Selken
// Current version: 	0.1
// File description:    AHB2APB bridge module global macros
// File history: 		0.1  - Dimitrije S. - Inital version.

	`define AHB_BUS_W  32
	`define AHB_ADDR_W 32
	`define APB_BUS_W  8
	`define APB_ADDR_W 32