// File name: 			AHB_Package.sv
// Creator name: 		Dimitrije Selken
// Current version: 	0.1
// File description:    AHB VIP module package
// File history: 		0.1  - Dimitrije S. - Inital version.

`ifndef AHB_PKG
`define AHB_PKG

`include "ahb_interface.sv"

package ahb_pkg;  

	import uvm_pkg::*;
	`include "uvm_macros.svh" 

	`include "ahb_transaction.sv"
	`include "ahb_master_driver.sv"
	`include "ahb_monitor.sv"
	`include "ahb_master_sequencer.sv"
	`include "ahb_master_agent.sv"

endpackage

`endif //ahb_pkg
